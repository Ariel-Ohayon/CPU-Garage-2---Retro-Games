library ieee;
use ieee.std_Logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_Logic_arith.all;

entity GAMEOVER is
port(
clk: in std_logic;
Xpxl,Ypxl: in std_logic_vector(31 downto 0);
topX,topY: in std_logic_vector(31 downto 0);
RGB: out std_logic_vector(11 downto 0);
drw: out std_logic);
end;

architecture one of GAMEOVER is
type mat is array (0 to 71, 0 to 301) of integer range 0 to 4095;
signal sRGB: mat :=
(
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,4095),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,0,0,0,0,0,0,0,0,0,0,0,0,0,0,4095),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,256,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,0,0,0,0,0,0,0,0,0,0,0,4095),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,0,0,0,0,0,0,0,0,0,0,4095),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,0,0,0,0,0,0,0,0,0,4095),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,0,0,0,0,0,0,0,0,4095),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,0,0,0,0,0,4095),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,512,512,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,0,0,0,0,4095),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,0,0,0,4095),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,0,0,0,4095),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,0,0,0,4095),
(0,0,0,0,0,0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,768,768,768,768,768,768,768,768,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,0,0,4095),
(0,0,0,0,0,0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,0,4095),
(0,0,0,0,0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,4095),
(0,0,0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,256,512,512,512,512,512,512,512,512,512,512,768,768,512,512,512,512,512,512,512,512,512,768,768,768,768,768,768,768,768,768,768,768,768,512,768,768,512,512,768,512,512,768,512,512,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,768,768,512,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,768,512,768,512,768,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,768,512,512,512,512,512,512,768,512,768,768,768,768,768,768,512,512,512,768,768,512,768,768,768,768,768,768,768,768,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,256,256,256,4095),
(0,0,0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,768,768,768,768,768,768,768,768,768,512,768,768,768,768,768,768,768,768,512,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,768,768,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,768,768,512,512,512,512,512,768,512,512,768,768,768,768,768,512,768,768,768,768,768,768,768,768,768,768,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,768,768,768,1024,768,1024,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,256,256,4095),
(0,0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,768,768,768,768,768,768,768,768,768,768,768,1024,768,768,1024,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,768,768,512,512,768,768,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,768,768,768,1024,768,768,1024,768,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,768,1024,1024,1024,1024,1024,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,768,768,512,512,512,512,512,512,512,512,512,512,512,512,256,512,256,256,256,256,256,256,256,256,256,256,4095),
(0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,768,512,512,512,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,769,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,768,768,768,768,768,768,768,768,768,768,768,1024,768,1024,768,768,768,768,768,768,768,768,768,768,1024,768,1024,768,1024,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,769,769,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,768,768,768,768,768,768,768,768,768,1025,1025,768,1024,1024,1024,1024,1024,768,1024,1024,768,1024,1024,768,1024,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,1024,1024,768,768,768,1024,1024,768,1024,1024,1024,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,4095),
(0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,513,769,512,512,768,768,768,768,512,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,769,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,768,1024,768,1024,768,1024,768,768,768,768,1024,1024,1024,1024,1024,1024,1024,768,1024,768,1024,768,1024,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,768,768,768,1024,768,1024,768,768,768,768,768,768,1024,768,768,768,768,768,768,768,768,768,1024,1024,1024,1024,768,768,768,1024,1024,1024,1024,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,768,768,1024,1024,1024,1024,768,1024,1024,1024,1024,768,768,1024,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,4095),
(0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,768,512,768,512,768,768,768,768,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,768,768,768,768,768,768,768,768,768,768,768,768,768,1025,769,768,768,768,1024,768,1024,1024,768,1024,1025,768,768,768,768,768,768,768,768,1024,1024,1025,768,1025,768,769,769,768,768,768,768,1024,768,1024,1024,1024,768,768,1025,768,768,768,1024,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,1024,1025,768,1025,768,769,769,768,768,768,768,1024,1024,768,1024,768,768,768,768,768,768,768,768,1024,768,768,768,1024,768,1024,1025,1024,1024,1024,768,1024,768,768,769,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,1024,1024,1024,768,1024,1024,1024,1024,768,1025,768,768,768,1024,1025,768,768,768,768,768,768,768,768,768,768,768,768,512,512,512,768,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,4095),
(0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,768,512,512,784,512,768,768,768,768,768,768,769,769,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,1024,1024,1024,1024,768,768,1024,768,768,768,1040,768,512,768,769,768,768,768,768,768,768,768,768,768,768,768,1024,768,768,1040,768,768,768,768,768,768,1024,1025,512,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,512,1024,768,768,768,768,768,768,1024,1040,768,1024,1025,1024,768,768,768,768,1040,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,512,768,769,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,1024,512,768,768,768,768,768,768,512,1040,768,768,1024,768,1024,1024,1024,1024,1024,768,512,1024,768,768,768,768,768,1024,768,768,768,768,768,1024,1024,1024,1024,1024,1024,1024,1024,769,768,1024,768,768,768,768,768,1024,768,768,768,1024,768,1024,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,1024,512,769,768,768,768,768,1040,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,768,768,769,513,768,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,4095),
(0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,784,2418,2691,3808,4064,4080,4080,4065,3792,2960,2144,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,768,768,1024,1024,768,1024,1569,4080,4080,4080,4066,2689,1040,768,769,1024,1024,1024,1024,1024,1024,1024,1024,768,768,768,768,768,1040,2674,2946,2688,2704,2704,2960,2704,2961,2417,1040,768,768,768,768,768,768,768,768,1024,768,768,1040,2417,2945,2704,2960,2704,2704,2960,2961,2673,1040,768,768,769,1025,768,768,1856,4051,4081,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4083,3506,1040,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1040,1842,2960,3248,3520,3520,3520,3520,3248,2976,2114,1040,768,768,768,1024,1024,768,768,768,768,1040,2417,2945,2688,2960,2960,2961,2690,1600,1024,768,768,768,768,768,768,768,768,768,768,768,768,1040,2674,2962,2944,2960,2960,2960,2945,768,1024,1025,768,1856,4050,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4080,4080,4080,4082,3506,1040,768,768,768,1024,1856,4051,4081,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4049,2960,1872,768,768,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,4095),
(0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,512,256,512,512,512,512,768,512,512,768,512,768,2688,4064,4080,4081,4080,4080,4080,4080,4080,4080,4080,4064,3792,2416,768,768,1024,1024,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,1024,768,768,2976,4080,4080,4081,4080,3808,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,768,768,4080,4080,4080,4080,4080,4080,4080,4080,4065,784,1024,768,768,1024,768,1024,1024,1024,1024,768,768,1328,4080,4064,4080,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,3520,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,769,768,768,769,768,2160,3792,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4064,2960,1312,769,1024,768,1026,1024,1024,768,1024,2688,4081,4080,4080,4080,4065,4080,2960,768,1024,1024,1024,1024,1024,1024,1024,768,768,1024,768,768,1600,4064,4080,4080,4080,4080,4080,3778,1024,768,768,768,1584,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4080,3776,768,1025,1024,768,768,1584,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,3248,1600,512,770,512,512,769,512,512,512,512,512,512,256,256,256,256,256,256,4095),
(0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,768,769,512,1872,3522,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4082,3506,1312,768,768,1024,768,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,768,1024,768,768,1040,3793,4080,4080,4080,4080,4080,2144,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,768,768,4080,4080,4080,4080,4080,4080,4080,4080,4082,2144,768,1024,768,1024,768,1024,1024,1024,1024,768,768,2145,4080,4080,4080,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4081,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4081,4080,3520,768,1024,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1312,3521,4080,4080,4081,4080,4081,4081,4080,4080,4081,4081,4080,4080,4064,4064,3794,2144,768,1024,768,1024,1024,768,768,1600,4081,4080,4080,4080,4080,4080,3520,768,1024,768,1024,768,768,768,768,1024,1024,1024,768,769,2688,4080,4080,4080,4080,4080,4080,2944,768,768,768,768,1584,4080,4080,4080,4080,4080,4081,4064,4080,4080,4081,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4080,3520,1024,1024,1024,768,768,1584,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,3521,1888,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,4095),
(0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,768,768,1872,3794,4080,4080,4080,4064,4080,4080,4080,4080,4080,4080,4080,4080,4065,4080,4080,4080,3794,1600,768,1025,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,768,2128,4082,4080,4080,4080,4080,4080,3505,768,768,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,768,768,4080,4080,4080,4080,4080,4080,4080,4080,4081,2976,768,768,1024,1024,768,1024,1024,1024,1024,768,768,3233,4080,4080,4080,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,3520,768,1024,1024,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,2128,4049,4064,4080,4080,4081,4080,4080,4080,4081,4081,4080,4080,4080,4080,4080,4080,4080,4064,2688,768,768,1024,1024,1024,768,768,3793,4064,4080,4080,4080,4081,4080,1312,768,768,1024,1024,1024,768,768,1024,1024,768,1024,768,3520,4080,4080,4080,4080,4080,4080,1584,768,1024,768,1024,1584,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4080,3520,768,768,1024,768,768,1584,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4064,4080,4081,4081,4080,4080,3793,1056,768,512,512,512,512,512,512,512,512,256,256,256,256,256,256,4095),
(0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,768,512,512,1600,4050,4080,4080,4064,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4064,4080,4080,3776,1312,768,768,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,768,768,1024,768,3248,4080,4080,4080,4080,4080,4080,4064,1312,768,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,768,768,4080,4080,4080,4080,4080,4080,4081,4080,4080,3792,1024,768,1025,768,1024,1024,1024,768,768,768,1040,3793,4080,4080,4080,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4064,4080,4080,4080,4080,4080,4080,4080,4080,4080,4064,4080,4081,3521,768,768,1024,768,768,768,768,768,768,768,768,1024,768,768,768,768,768,768,1024,768,1584,3776,4080,4080,3808,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4064,4080,4080,2400,769,768,768,768,1024,768,2960,4080,4080,4080,4080,4080,4080,2416,768,1024,1024,1024,1024,1024,768,768,768,768,768,1312,4080,4080,4080,4080,4080,4080,3792,1024,769,1024,768,1024,1584,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,3520,768,768,1024,768,768,1584,4080,4080,4080,4080,4081,4064,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4064,4080,4080,2976,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,4095),
(0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,256,512,512,768,3520,4080,4080,4080,4080,4080,4080,4064,4080,4080,4080,4064,4081,4081,4064,4080,4080,4081,4081,4080,4080,3233,768,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,768,768,1312,4064,4080,4080,4080,4080,4080,4080,4080,2688,768,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,768,768,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,1584,768,1025,768,1024,1024,1024,768,768,1024,1856,4080,4080,4080,4081,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4080,4080,3792,4082,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4065,3504,1040,1024,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,1024,768,768,3249,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4064,4080,4050,1312,768,768,768,1024,768,1584,4080,4080,4080,4080,4080,4080,3520,768,1024,1024,768,768,1024,768,768,1024,768,768,2416,4080,4080,4080,4080,4080,4080,2688,768,769,1024,1024,1024,1584,4080,4080,4080,4064,4080,4080,4080,4048,4065,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4081,3232,1040,768,1024,768,768,1584,4080,4080,4080,4080,4064,4080,4080,4064,4081,4080,4080,4080,4080,4080,4080,4064,4080,4080,4080,4080,4080,4080,4080,4081,1328,512,768,512,512,512,512,512,512,512,512,256,256,256,256,4095),
(0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,768,2416,4080,4080,4064,4080,4080,4064,4080,4080,4080,4080,4081,4081,4064,4080,4080,4080,4080,4064,4080,4080,4080,4064,2400,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,768,2672,4080,4080,4080,4080,4064,4080,4080,4080,3520,768,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,768,768,4080,4080,4080,4080,4080,4064,4080,4080,4080,4080,2688,768,768,768,768,768,768,768,768,1024,2688,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4064,2976,1040,768,768,768,768,768,768,768,768,768,768,768,768,1024,768,1024,1040,768,1024,1024,768,768,768,768,768,768,768,768,768,768,768,768,1024,1024,768,768,2144,4081,4080,4064,4080,4080,4080,4080,4080,4080,4080,3792,3776,4064,4081,4065,4080,4080,4064,4080,4080,4080,4080,2976,768,768,1024,1024,1024,768,3792,4080,4080,4080,4080,4080,4080,1312,768,1024,1024,768,1024,1024,1024,1024,768,1024,3520,4080,4080,4080,4080,4080,4081,1600,768,1024,1024,1024,768,1584,4080,4080,4080,4080,4080,4065,3233,1040,768,768,768,768,768,768,768,768,768,768,1025,768,768,768,768,1040,768,1025,1024,768,768,1584,4080,4080,4080,4080,4080,4065,2976,1040,768,768,768,769,1024,768,769,1040,2432,4081,4080,4080,4080,4080,4080,4080,2960,512,513,512,512,512,512,512,512,512,512,512,256,256,256,4095),
(0,0,0,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,784,3520,4080,4080,4081,4080,4080,4080,4080,4080,2960,1584,768,768,1312,2960,4065,4080,4080,4080,4080,4080,4080,4080,3521,768,1024,1024,1024,1024,1024,1024,1024,1024,768,768,1024,768,1024,3776,4080,4080,4080,4080,4080,4080,4080,4080,4064,1600,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,768,768,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,3777,768,768,768,768,768,768,1024,768,768,3776,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4080,3232,768,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,768,768,1025,1024,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,768,768,1024,3536,4080,4080,4080,4081,4064,4080,4064,4049,2416,1040,768,768,768,2128,3504,4080,4080,4081,4080,4080,4080,4080,4080,1328,768,1024,1024,1024,768,2689,4080,4080,4080,4080,4080,4080,2672,768,1024,1024,768,1024,768,1024,768,768,1568,4080,4081,4080,4080,4081,4080,3777,1040,768,768,1024,768,768,1584,4080,4080,4080,4080,4080,4080,3232,768,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,768,1024,1024,1024,768,768,1584,4080,4080,4080,4080,4080,4080,3233,768,768,768,1024,768,768,1024,1025,768,1056,2688,4065,4080,4064,4080,4064,4080,3520,768,512,768,512,512,512,512,512,512,512,512,256,256,256,4095),
(0,0,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,769,1600,4080,4066,4080,4080,4080,4080,4080,3793,1600,768,768,768,769,769,768,1856,3778,4080,4080,4080,4080,4064,4080,4065,1872,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1841,4064,4080,4080,4080,4080,4080,4081,4080,4080,4081,2688,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,768,768,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4065,768,768,1024,1024,1024,768,768,1024,768,4081,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4081,4081,3232,768,769,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1025,768,1025,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,768,768,1024,768,768,1024,1569,4080,4080,4080,4080,4080,4080,4064,3792,1312,1024,768,768,1025,768,768,1024,3248,4080,4080,4080,4080,4080,4080,4080,2417,768,1024,1024,768,1024,1584,4080,4080,4080,4080,4080,4080,3505,768,1024,768,768,768,768,1024,768,1024,2402,4080,4081,4080,4080,4080,4064,2961,768,768,768,1024,768,768,1856,4080,4080,4080,4080,4080,4080,3232,768,769,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,768,768,1024,768,1024,768,768,1584,4080,4080,4080,4080,4080,4080,3232,768,768,768,768,1024,1024,1024,768,1024,768,1584,4066,4080,4080,4080,4080,4080,4081,1056,768,512,512,512,512,512,512,512,512,512,256,256,256,4095),
(0,0,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,2976,4080,4080,4080,4080,4080,4080,4066,1584,768,768,1024,1024,768,1024,768,768,1584,3808,4081,4080,4080,4080,4081,4065,2720,768,1024,1024,768,1024,1024,1024,1024,1024,1024,768,768,2976,4080,4080,4080,4080,4081,4080,4080,4080,4081,4080,3808,768,768,768,1024,768,1024,768,1025,768,1024,1024,1024,768,768,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,2144,768,1024,1024,1024,768,1024,768,2416,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4080,3248,768,768,768,1024,768,768,768,768,768,768,768,768,1024,1025,1024,1024,768,1024,768,768,1024,1024,1024,1024,1024,1024,1024,1024,768,768,1024,1024,768,1024,768,2960,4080,4080,4080,4080,4080,4080,4050,1312,1024,1024,1024,1024,1024,1024,1024,1024,1024,3506,4080,4080,4080,4080,4080,4080,3504,768,1024,768,1024,768,1024,3777,4080,4081,4080,4081,4080,4064,1024,768,768,1024,1024,1024,768,1024,768,3248,4080,4080,4080,4081,4080,4081,1312,1024,1024,1024,1024,1024,768,1584,4080,4080,4080,4080,4080,4080,3233,1024,1024,1024,768,768,768,768,768,768,768,768,1024,1024,1025,768,1025,768,768,768,1024,768,768,1584,4080,4080,4080,4080,4080,4080,3233,768,1024,1024,1024,768,1024,1024,768,1024,1024,768,3520,4080,4080,4080,4064,4080,4080,1872,768,768,512,512,512,512,512,512,512,512,256,256,256,4095),
(0,0,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,3232,4080,4080,4080,4080,4080,4080,3248,1040,768,1024,768,1024,768,768,768,768,1024,3248,4064,4080,4080,4080,4081,4081,3520,768,1024,1024,1024,1024,768,768,1024,768,768,768,784,3793,4080,4064,4080,4080,4080,4080,4080,4080,4080,4080,4080,2145,768,1025,1024,1024,1024,768,768,768,1024,1024,1024,768,768,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,2960,768,1024,768,1024,768,1024,768,3232,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4080,3232,768,1025,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,768,768,1024,768,768,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,768,768,768,3232,4080,4080,4080,4080,4080,4080,2976,768,1024,1024,1024,1024,1024,1024,1024,1024,768,2416,4080,4080,4080,4080,4080,4080,3792,768,1024,768,1024,768,768,2944,4080,4080,4080,4080,4080,4080,2401,1024,768,1024,768,768,1024,768,1040,3792,4080,4080,4080,4080,4080,3520,1040,768,1024,1024,1024,1024,768,1584,4080,4080,4080,4080,4080,4080,3232,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,768,1024,1024,768,1024,768,768,1584,4080,4080,4080,4080,4080,4080,3233,768,1024,768,1024,1024,1024,768,1025,1024,768,768,3232,4064,4080,4080,4080,4080,4080,2144,512,768,512,512,512,512,512,512,512,512,256,256,256,4095),
(0,0,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,768,3520,4080,4080,4080,4080,4080,4064,2416,768,768,1024,1024,1024,768,768,1024,768,768,768,1024,1024,768,768,768,1024,768,1024,1024,768,1024,1024,768,768,1024,1024,768,768,2144,4081,4080,4080,4080,4080,4080,3792,4080,4080,4080,4081,4080,3233,768,768,768,1024,1024,768,768,768,1024,1024,1024,768,768,4080,4080,4080,4080,4080,4080,4065,4080,4080,4080,4080,3792,768,1024,1024,1024,1024,768,768,4048,4065,4080,4080,4080,3792,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4080,3232,768,769,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1025,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,768,768,768,3504,4080,4080,4080,4080,4080,4080,2144,768,1024,1024,1024,1024,1024,1024,1024,1024,768,1040,4064,4080,4080,4080,4080,4080,4080,768,768,1024,768,1024,768,1584,4080,4080,4080,4080,4080,4080,3232,768,1024,768,1024,768,1024,768,2144,4080,4080,4080,4080,4080,4080,2688,1024,768,1024,1024,1024,1024,768,1584,4080,4080,4080,4080,4080,4080,3232,768,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,768,768,768,768,1024,768,768,1584,4080,4080,4080,4080,4080,4080,3232,1024,1024,768,1024,768,768,1024,1024,1024,1024,768,3232,4080,4080,4080,4080,4080,4080,2145,512,768,512,512,512,512,512,512,512,512,256,256,256,4095),
(0,0,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,768,3792,4080,4080,4080,4080,4080,4081,1856,768,1024,1024,1024,1024,768,1024,1024,1024,1024,1024,1024,768,768,1024,1024,768,1024,1024,768,768,768,768,1024,1024,1024,1024,768,768,3504,4080,4080,4081,4080,4080,3792,2704,4080,4080,4080,4080,4080,4065,1312,768,768,1024,768,768,768,768,1024,1024,1024,768,768,4080,4080,4080,4080,4080,4080,3249,4080,4080,4080,4080,4080,1584,768,1024,768,768,768,1600,4080,4064,4080,4080,4080,2704,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4081,4080,4080,3232,768,1025,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,768,768,768,1024,1025,768,768,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,768,768,768,3521,4080,4080,4080,4080,4080,4081,1584,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,512,3792,4080,4080,4080,4081,4080,4080,768,768,1024,768,1024,769,1024,3792,4080,4080,4080,4080,4064,4064,1040,1025,768,1024,1024,768,768,3504,4080,4080,4080,4080,4080,4080,1600,768,1025,1024,1024,768,1024,768,1584,4080,4080,4080,4080,4080,4080,3232,768,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,768,1024,768,1024,1024,1024,1024,768,768,1584,4080,4080,4080,4080,4080,4080,3232,768,768,768,768,769,1025,1024,768,1024,768,1024,3520,4080,4080,4080,4080,4080,4081,1856,512,768,512,512,512,512,512,512,512,512,256,256,256,4095),
(0,0,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,3792,4080,4081,4080,4080,4080,4081,1584,768,768,1024,1024,1024,768,1024,1024,1024,768,768,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,768,768,768,768,768,768,768,1312,4064,4080,4080,4080,4080,4080,2688,1328,4080,4080,4080,4080,4080,4080,2689,768,1024,1024,768,768,1024,768,1024,1024,1024,768,768,4080,4080,4080,4080,4080,4080,2144,4081,4080,4080,4081,4080,2688,768,1024,768,1024,1024,2688,4080,4080,4080,4081,4080,1600,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4080,3232,768,768,1024,1024,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,768,768,768,3520,4080,4080,4080,4080,4064,4081,1024,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,769,3520,4080,4080,4080,4080,4080,4080,768,768,1024,768,1024,1025,768,2688,4080,4064,4080,4080,4080,4080,2400,1025,768,768,1024,768,768,4065,4080,4080,4081,4080,4080,3520,1024,768,768,1024,1024,768,1024,768,1584,4080,4080,4064,4080,4080,4081,3232,768,768,1024,768,768,768,768,768,768,768,768,768,768,768,1024,1024,1024,768,768,1024,768,768,1584,4080,4080,4080,4080,4080,4080,3232,768,1024,768,768,768,1024,1024,1024,1025,512,1312,4065,4080,4080,4080,4080,4080,4082,1312,512,768,512,512,512,512,512,512,512,512,256,256,256,4095),
(0,0,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,3792,4080,4080,4080,4080,4080,4081,1584,1024,768,768,768,1024,1024,768,768,1025,768,768,1024,1024,768,768,768,768,768,768,768,1024,1024,768,768,1024,768,1024,768,2689,4080,4080,4080,4080,4080,4064,1584,512,3777,4080,4080,4080,4080,4080,3521,768,768,768,1024,1024,1024,768,1024,1024,1024,768,768,4080,4080,4080,4080,4081,4080,1056,4065,4080,4080,4080,4080,3504,768,768,1025,1024,768,3520,4064,4080,4064,4080,3792,768,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4065,3232,1040,768,768,768,768,768,768,768,768,768,768,768,768,1040,512,768,768,1024,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,768,1024,1024,768,768,3520,4080,4080,4080,4080,4080,4080,768,768,1024,1024,1024,1024,1024,1024,1024,1024,768,1025,3504,4080,4080,4080,4080,4080,4064,768,1024,1024,1024,1024,1024,768,1600,4081,4080,4080,4080,4080,4080,3248,768,1024,1024,1024,1024,1856,4080,4080,4080,4081,4080,4080,2688,768,1024,768,1024,1024,1024,1024,768,1584,4080,4080,4080,4080,4080,4065,2960,1040,768,768,768,768,768,768,768,768,768,768,768,768,1040,768,1026,768,768,1024,1024,768,768,1584,4080,4080,4080,4080,4080,4080,3233,768,768,1025,768,768,768,768,1025,768,1296,2688,4080,4080,4080,4080,4080,4080,3794,768,768,512,512,512,512,512,512,512,512,512,256,256,256,4095),
(0,0,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,3792,4080,4080,4080,4080,4080,4080,1584,1024,768,768,768,768,768,1040,768,768,768,768,768,768,768,768,768,768,768,1024,768,768,1024,1024,1024,1024,1024,768,1040,3776,4080,4080,4080,4080,4080,3520,1024,768,2416,4080,4080,4080,4080,4080,4080,1872,768,768,1024,1024,1024,768,1024,1024,1024,768,768,4080,4080,4080,4080,4081,4080,768,3248,4080,4080,4080,4080,3792,1040,768,1024,768,1024,4080,4080,4080,4080,4080,2960,768,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4080,4080,4065,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4050,1040,768,768,1024,1024,1025,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,1024,768,768,3520,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,768,3520,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,1024,1024,768,768,3520,4080,4080,4080,4080,4080,3792,1024,768,1024,768,1024,2976,4080,4080,4080,4080,4080,4064,1600,768,1024,1024,1024,1024,1024,1024,768,1584,4080,4080,4081,4080,4080,4080,4080,4065,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4080,4049,1040,768,1024,1024,768,1024,768,768,1584,4080,4080,4080,4080,4080,4080,3232,1040,768,768,768,768,768,768,768,1040,2689,4066,4080,4080,4080,4080,4080,4080,2704,512,768,768,512,512,512,512,512,512,512,512,256,256,256,4095),
(0,0,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,768,512,3792,4080,4080,4080,4080,4080,4080,1584,768,768,768,768,768,1856,4050,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,1570,1024,768,1024,1024,1024,768,768,768,1857,4064,4080,4065,4081,4080,4080,2960,768,769,1312,4080,4080,4080,4080,4080,4080,2960,1025,768,1024,769,1024,768,1024,1024,1024,768,768,4080,4080,4080,4080,4065,4080,768,2704,4080,4081,4080,4080,4080,2128,1024,768,1024,2401,4080,4080,4080,4080,4080,1872,768,4065,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4080,4080,4082,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,768,768,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,768,768,768,3520,4080,4080,4080,4080,4080,4080,1025,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,768,3776,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,1024,1024,768,768,2960,4080,4080,4081,4080,4080,4080,2113,768,1024,768,1024,3792,4080,4080,4080,4080,4080,3792,768,768,768,1024,1024,1024,1024,1024,768,1584,4080,4080,4080,4080,4080,4080,4080,4065,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4082,768,768,768,1024,1024,1024,768,768,1584,4080,4080,4080,4080,4081,4080,4080,4049,4080,4080,4080,4080,4080,4064,4080,4081,4080,4080,4080,4081,4080,4080,4080,4080,1872,512,768,768,512,512,512,512,512,512,512,512,256,256,256,4095),
(0,0,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,768,3808,4080,4080,4080,4080,4080,4080,1584,768,768,1024,1024,768,1584,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,1600,768,1024,1024,1025,1024,1024,1024,768,3232,4080,4064,4065,4081,4080,4080,1312,768,768,768,3520,4064,4080,4081,4081,4080,4064,784,768,768,1024,1024,768,1024,1024,1024,768,768,4080,4080,4080,4080,4081,4080,768,1312,4081,4080,4080,4080,4080,2976,768,768,768,3232,4080,4080,4080,4065,4064,1024,768,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,768,768,768,1024,768,768,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,1024,768,768,3520,4080,4064,4080,4080,4080,4080,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,3520,4080,4080,4080,4080,4080,4080,768,768,1024,1024,1024,768,768,1024,1312,4081,4080,4081,4080,4080,4080,3232,768,768,768,1872,4080,4080,4080,4080,4080,4081,2944,768,768,1024,768,1024,1024,1024,1024,768,1584,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,768,768,1024,1024,1024,1024,768,768,1584,4080,4080,4080,4080,4080,4080,4064,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4080,4080,4080,2976,784,512,768,768,512,512,512,512,512,512,512,512,256,256,256,4095),
(0,0,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,768,3808,4080,4080,4080,4080,4080,4080,1584,768,1024,1024,1024,768,1584,4080,4080,4081,4081,4080,4081,4081,4080,4064,4080,4080,4080,1584,768,768,1024,1024,768,1024,1024,768,4064,4080,4081,4080,4080,4080,3520,1024,768,768,1024,2688,4080,4080,4080,4081,4080,4081,2144,768,1024,1024,1024,768,1024,1024,1024,768,768,4080,4080,4080,4080,4080,4080,768,1024,3504,4080,4080,4080,4080,3776,1024,768,768,3792,4080,4080,4080,4081,3504,1024,768,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4064,4080,768,768,1024,768,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,1024,768,768,3520,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,3520,4080,4080,4080,4080,4080,4080,768,768,1024,1024,1024,768,768,768,1040,3520,4080,4080,4080,4080,4080,3792,1024,768,768,2960,4080,4080,4080,4080,4080,4064,1856,768,768,768,768,1024,1024,1024,1024,768,1584,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,768,1025,768,768,1024,1024,768,768,1584,4080,4080,4080,4080,4064,4080,4080,4080,4081,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4064,4080,3521,1328,512,768,512,768,512,512,512,512,512,512,512,512,256,256,256,4095),
(0,0,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,768,3808,4080,4080,4080,4080,4080,4080,1584,768,1024,768,768,768,1584,4081,4080,4080,4080,4080,4080,4080,4081,4080,4080,4080,4080,1584,768,768,1024,1024,1024,1025,1024,2144,4082,4080,4081,4080,4080,4080,2688,768,768,768,768,1312,4064,4080,4080,4080,4080,4080,3505,768,768,768,1024,768,1024,1024,1024,768,768,4080,4080,4080,4080,4080,4080,768,1024,2688,4080,4080,4080,4080,4080,1584,768,1584,4080,4080,4080,4080,4080,2144,768,768,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,768,768,1025,1024,768,768,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,1024,768,768,3520,4064,4080,4080,4080,4080,4080,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,3520,4080,4080,4080,4080,4080,4080,768,768,1024,1024,1024,768,768,768,1024,2688,4080,4080,4080,4080,4080,4081,1856,768,768,4048,4080,4080,4081,4080,4080,3792,1024,1024,1024,768,1024,1024,1024,1024,1024,768,1584,4080,4080,4081,4080,4080,4080,4080,4081,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4081,768,769,1024,1024,1024,1024,768,768,1584,4080,4080,4080,4080,4081,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,3777,1873,768,512,768,768,768,512,512,512,512,512,512,512,512,256,256,256,4095),
(0,0,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,768,3792,4080,4080,4080,4080,4080,4080,1584,768,1024,1024,1024,768,1584,4081,4080,4080,4080,4080,4080,4080,4081,4080,4080,4080,4081,1584,768,1024,1024,768,1024,769,768,3520,4064,4080,4080,4081,4080,4064,1312,768,1024,1024,1024,768,3505,4080,4080,4080,4080,4080,4064,1328,768,1024,1024,768,1024,1024,1024,768,768,4080,4080,4080,4080,4080,4080,768,768,1584,4080,4080,4080,4080,4080,2416,768,2689,4080,4080,4080,4080,4064,1296,768,768,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4080,4080,4064,4081,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4064,1040,768,1024,768,768,768,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,1024,768,768,3520,4080,4080,4080,4080,4080,4064,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,3520,4080,4080,4080,4080,4080,4080,768,768,1024,1024,1024,768,768,1025,768,1600,4080,4080,4080,4080,4080,4080,2960,768,1584,4080,4080,4080,4080,4080,4080,2704,768,1024,1024,1024,1024,1024,1024,768,1024,768,1584,4080,4080,4081,4080,4080,4080,4080,4064,4081,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4048,1040,768,1024,1024,768,1024,768,768,1584,4080,4080,4080,4080,4080,4064,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4065,4065,3248,1328,768,768,768,768,512,768,512,512,512,512,512,512,512,512,256,256,256,4095),
(0,0,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,3792,4080,4080,4080,4080,4080,4080,1584,768,1024,768,768,768,1600,4049,4081,4080,4080,4066,4080,4080,4080,4080,4080,4080,4081,1584,768,1024,768,768,1024,768,1568,4080,4080,4080,4080,4064,4080,3520,768,1024,768,768,1024,1024,2416,4080,4080,4080,4080,4080,4080,2688,768,1024,1024,768,1024,1024,1024,768,768,4080,4080,4080,4080,4080,4080,768,768,1024,3520,4081,4080,4080,4080,3248,512,3505,4080,4080,4080,4080,3520,768,1024,768,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4081,3233,1040,768,768,1025,768,768,768,768,768,768,768,768,768,1040,512,1024,1024,1024,768,768,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,1024,768,768,3520,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,3520,4080,4080,4080,4080,4080,4080,768,768,1024,1024,1024,768,768,768,768,1024,3520,4080,4080,4081,4080,4080,3793,768,2688,4080,4080,4080,4080,4080,4064,1584,1024,768,768,1024,768,1024,1024,768,1024,768,1584,4080,4080,4080,4080,4080,4064,3233,1040,768,768,768,768,768,768,768,768,768,768,768,768,1040,769,769,1024,768,1024,1024,768,768,1584,4080,4080,4080,4080,4080,4080,4080,4064,4080,4081,4065,4080,4080,4080,4080,4080,4080,4064,3248,1872,1040,768,512,768,768,512,768,512,512,512,512,512,512,512,512,512,256,256,256,4095),
(0,0,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,3792,4080,4080,4080,4080,4080,4080,1584,768,768,1024,768,768,512,1040,768,768,768,1040,3248,4080,4082,4080,4080,4080,4080,1584,768,1024,1024,1024,768,768,2688,4081,4080,4080,4080,4080,4080,2416,768,768,768,1024,1025,768,1312,3808,4080,4080,4080,4080,4080,3792,768,768,768,768,1024,1024,1024,768,768,4080,4080,4080,4080,4080,4080,1024,1024,1024,2689,4081,4080,4081,4080,4064,1040,4064,4080,4080,4080,4080,2689,768,1024,768,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4080,3232,768,768,1024,768,768,768,768,768,768,768,768,768,768,768,1025,1024,768,768,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,1024,768,768,3520,4080,4080,4080,4080,4080,4080,768,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,3520,4080,4080,4080,4080,4080,4080,768,768,1024,1024,1024,768,768,768,1024,768,2688,4080,4080,4081,4080,4080,4080,1584,3792,4080,4080,4080,4080,4080,3793,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,1584,4080,4080,4080,4080,4080,4080,3233,768,768,1024,768,768,768,768,768,768,768,768,1024,768,768,1024,768,768,768,1024,1024,768,768,1584,4080,4080,4080,4080,4080,4080,3234,1024,768,768,1600,4081,4080,4080,4080,4080,4080,4080,3248,784,768,768,1024,768,768,768,512,768,512,512,512,512,512,512,512,512,256,256,256,4095),
(0,0,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,3792,4080,4080,4080,4080,4080,4080,1600,768,768,1024,1024,768,768,768,768,1024,1024,768,3777,4080,4064,4080,4080,4080,4080,1584,768,1024,1024,768,768,1040,3520,4080,4080,4080,4081,4080,3792,1584,768,768,1024,1024,768,768,1040,3233,4066,4080,4080,4080,4080,4080,1872,768,1024,768,1024,1024,1024,768,768,4080,4080,4080,4080,4080,4080,768,1024,768,1584,4080,4080,4080,4080,4080,2688,4080,4080,4080,4080,3808,1584,1024,1024,768,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4080,3248,768,768,1024,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,1024,768,768,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,1024,768,768,3520,4080,4080,4080,4080,4080,4080,1296,768,1024,1024,1024,1024,1024,1024,1024,1024,768,768,3792,4080,4080,4080,4080,4080,4080,768,768,1024,1024,1024,768,768,1024,1024,768,1600,4064,4080,4080,4080,4080,4080,2976,4080,4081,4080,4080,4080,4080,2689,768,768,1024,1024,1024,1024,1024,1024,1024,1024,768,1584,4080,4080,4080,4080,4080,4080,3232,768,769,768,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,768,1024,1024,1024,1024,768,768,1584,4080,4080,4080,4080,4080,4080,3233,768,1024,768,1024,2688,4081,4080,4080,4080,4080,4080,4065,2416,1025,768,768,768,768,512,769,768,512,512,512,512,512,512,512,512,256,256,256,4095),
(0,0,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,3792,4080,4080,4080,4080,4080,4081,1600,1024,768,1024,1024,1024,1025,768,1025,1024,1024,768,4050,4080,4080,4080,4080,4080,4080,1312,768,1024,1024,768,1024,1856,4080,4080,4081,4080,4064,4080,4080,4066,4065,4081,4080,4064,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,2960,1025,768,768,1024,1024,1024,768,768,4080,4080,4080,4080,4080,4080,768,1024,1024,768,3808,4080,4080,4080,4080,4081,4080,4080,4080,4080,3536,512,1024,768,768,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4080,3232,768,769,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,768,1024,768,768,768,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,1024,768,768,3520,4080,4080,4080,4080,4080,4080,1858,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,3792,4080,4080,4080,4080,4080,4080,768,768,1024,1024,1024,768,768,1024,768,768,768,3792,4080,4080,4080,4080,4081,4080,4080,4064,4080,4080,4080,4080,1584,768,768,1024,1024,1024,768,1024,1024,1024,1024,768,1584,4080,4080,4080,4080,4080,4080,3249,768,1025,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1025,768,1024,1024,768,768,1024,768,768,1584,4080,4080,4080,4080,4080,4080,3234,1024,768,1024,769,1312,3808,4080,4080,4081,4081,4080,4080,3793,768,1024,768,768,769,768,768,512,512,512,512,512,512,512,512,512,256,256,256,4095),
(0,0,0,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,513,768,3248,4080,4080,4080,4064,4080,4080,2688,768,769,768,1024,768,1024,1024,1024,768,1024,2416,4080,4080,4080,4080,4080,4081,4064,768,1025,1024,1024,1024,768,2976,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4080,4080,4082,4080,4064,768,768,768,768,768,1024,768,769,4080,4080,4080,4080,4080,4080,768,768,1024,1024,2976,4080,4080,4065,4081,4080,4080,4080,4080,4080,2688,1024,768,768,768,4064,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4080,3248,768,1025,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,768,768,768,768,768,768,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,3505,4080,4080,4081,4081,4080,4080,2689,768,768,768,1024,1024,768,768,768,1024,768,1584,4064,4080,4064,4080,4080,4080,4081,768,768,1024,768,768,1024,768,768,1024,768,768,2944,4081,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,3778,768,768,768,768,768,768,1024,1024,1024,1024,1024,768,1584,4080,4080,4080,4080,4080,4080,3232,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,768,1024,1024,768,1024,768,1024,768,768,1584,4080,4080,4080,4080,4080,4080,3232,768,768,1024,1024,1024,2417,4081,4080,4080,4080,4080,4080,4064,2960,512,768,768,768,768,512,768,512,512,512,512,512,512,512,512,256,256,256,4095),
(0,0,0,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,768,2960,4080,4064,4080,4081,4064,4080,3793,1328,768,1024,768,1025,1025,768,1024,768,1024,3520,4081,4080,4064,4080,4080,4081,3792,1024,768,1024,1024,768,768,3793,4080,4080,4080,4080,4080,4080,4080,4081,4081,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4080,4080,2144,768,768,768,768,1024,768,768,4080,4080,4080,4080,4080,4080,768,768,1024,1024,1872,4080,4080,4080,4080,4080,4080,4081,4080,4064,1584,768,1024,1024,768,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4080,3248,768,1024,768,1024,768,768,768,768,768,768,768,768,1024,768,768,1024,768,768,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,768,768,768,2960,4080,4080,4080,4080,4080,4080,3504,1040,1024,1024,1024,1024,1024,1024,768,768,768,2960,4080,4080,4080,4080,4080,4080,3776,768,768,768,768,768,768,768,768,768,768,768,1856,4064,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,2945,768,768,768,768,768,768,1024,1024,1024,1024,1024,768,1584,4080,4080,4080,4080,4080,4080,3248,768,768,768,768,768,768,768,768,768,768,768,1024,1024,768,768,1024,768,768,768,1024,768,768,1584,4080,4080,4080,4080,4080,4080,3232,768,768,1024,1024,1024,1040,3521,4080,4080,4080,4080,4080,4080,4066,1856,768,768,768,512,768,768,512,512,512,512,512,512,512,512,256,256,256,4095),
(0,0,0,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,768,2144,4081,4080,4080,4080,4080,4080,4081,3248,1584,768,768,768,768,768,768,1040,3234,4080,4080,4080,4080,4081,4080,4081,2704,1024,1024,1024,1024,1025,2144,4082,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,3505,768,1024,768,768,1024,768,768,4080,4080,4080,4080,4080,4080,768,768,1024,1024,768,4065,4080,4080,4080,4080,4080,4080,4080,3793,768,769,1024,1024,768,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4080,3232,768,1024,768,768,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,768,1024,1024,1024,768,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,2400,4080,4064,4080,4080,4080,4080,4081,2688,1024,768,768,768,1024,1024,768,768,1872,4064,4080,4080,4080,4080,4080,4080,2960,1024,768,768,1024,768,1024,768,1024,768,1024,1024,1024,3792,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,1584,768,768,768,1024,768,768,1024,1024,1024,1024,1024,768,1584,4080,4080,4080,4080,4080,4080,3233,768,768,1025,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,1024,768,1024,1024,1024,768,768,1584,4080,4080,4080,4080,4080,4080,3232,768,768,1024,1024,1024,768,2144,4081,4080,4080,4080,4064,4081,4080,3232,768,768,512,768,768,768,512,512,512,512,512,512,512,512,256,256,256,4095),
(0,0,0,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,1328,3794,4064,4081,4064,4080,4080,4080,4080,3793,2946,1312,768,768,1040,2689,3793,4064,4080,4080,4080,4080,4064,4080,4081,1584,1024,1024,768,768,768,3520,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4064,4080,4080,4080,4080,4065,1312,768,1024,768,768,1024,768,4080,4080,4080,4080,4080,4080,768,768,1024,1024,512,3248,4080,4080,4080,4081,4080,4080,4080,3233,769,1025,768,768,768,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4081,3232,768,768,768,1026,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,768,768,1024,1024,768,768,768,768,768,768,768,768,768,1024,1024,768,768,768,768,768,1040,4064,4080,4080,4080,4080,4080,4081,4080,2672,1056,512,769,769,512,1040,2144,4065,4080,4080,4080,4080,4080,4064,4080,2128,1024,768,768,1024,1024,1024,1024,1024,1024,1024,1024,768,2704,4080,4080,4080,4080,4080,4080,4080,4080,4080,3793,1024,768,1024,768,1024,768,1024,1024,1024,1024,768,1024,768,1584,4080,4080,4080,4080,4080,4080,2976,768,768,1025,1024,1024,1024,1024,1024,1024,1024,1024,768,768,1024,1025,768,768,1024,1024,1024,768,768,1584,4080,4080,4080,4080,4080,4080,3232,768,768,1024,1024,1024,768,1024,3249,4080,4080,4080,4080,4080,4080,4080,2416,513,768,768,768,512,512,512,512,512,512,512,512,512,256,256,256,4095),
(0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,768,2688,4080,4080,4080,4080,4081,4080,4064,4080,4081,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,3232,768,1024,768,1024,768,1312,4080,4080,4080,4081,4080,4080,4081,4064,4081,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4065,4081,4080,4080,4080,4080,4080,2688,768,768,1024,768,1024,768,4080,4080,4080,4080,4080,4080,768,768,1024,1024,1040,2144,4080,4080,4080,4080,4080,4081,4080,1856,1024,1024,768,768,768,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4064,2976,1040,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,1024,512,1025,1024,768,768,768,768,768,768,768,768,1024,1024,768,1024,768,1024,1024,768,2704,4080,4080,4064,4080,4080,4064,4080,4081,3792,2960,2144,2144,2960,3504,4065,4080,4080,4080,4080,4080,4080,4080,3792,1024,768,768,768,1024,768,768,1024,768,1024,768,768,1024,1584,4064,4080,4080,4080,4080,4080,4080,4080,4081,2704,768,768,1024,768,1024,768,1024,1024,1024,1024,768,1024,768,1584,4080,4080,4080,4080,4081,4081,2976,1040,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,1040,768,1024,1024,768,768,1584,4080,4080,4080,4080,4080,4080,3232,768,768,1024,1024,1024,768,768,1584,4064,4080,4080,4080,4080,4080,4080,3792,768,768,512,768,512,512,512,512,512,512,512,512,256,256,256,256,4095),
(0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,768,512,1312,3808,4080,4080,4080,4064,4081,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4064,4080,4066,1584,768,1024,1024,1024,768,2688,4080,4080,4080,4080,4080,4065,2961,1040,768,768,768,768,768,768,768,768,768,768,768,2128,4081,4080,4080,4080,4080,4080,3793,1024,768,1024,1024,1024,768,4080,4080,4080,4080,4080,4080,768,768,1024,1024,769,1024,3793,4080,4080,4080,4080,4080,4065,768,768,1024,1024,768,768,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4081,4080,4080,4080,3792,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4065,4064,3505,1040,768,768,1024,1024,1024,1024,1024,1024,1024,1024,768,768,768,768,768,1024,1024,768,1312,4064,4080,4065,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4080,4080,4080,4080,4080,4080,4080,2144,768,768,1024,1024,768,768,768,1024,1024,1024,1024,1024,1024,1024,3793,4080,4080,4080,4080,4080,4064,4080,4066,1600,768,768,1024,1024,1024,768,1024,1024,1024,1024,1024,1024,768,1584,4080,4080,4065,4080,4080,4080,4080,4064,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4064,3504,1040,768,1024,768,768,1584,4080,4080,4080,4080,4080,4080,3232,768,768,1024,1024,1024,1024,1025,768,2704,4080,4080,4080,4080,4080,4080,4080,2688,512,768,768,768,512,512,512,512,512,512,256,256,256,256,256,4095),
(0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,513,512,512,2144,4066,4080,4080,4080,4080,4080,4081,4080,4081,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4065,2689,1024,768,1024,1024,768,784,3792,4080,4080,4080,4080,4080,4082,2128,768,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,3793,4080,4080,4080,4080,4080,4080,1856,768,1024,1024,768,768,4080,4080,4080,4080,4080,4080,768,768,1024,1024,768,1040,3232,4064,4081,4080,4080,4064,2961,1024,1024,1024,1024,768,768,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4080,4080,4065,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4080,3778,768,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,768,768,768,768,768,1024,1025,768,2688,4064,4081,4064,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,3232,768,1024,1024,1024,1024,768,1024,1024,1024,1024,1024,1024,1024,768,768,2689,4080,4080,4080,4080,4080,4080,4080,3521,768,1024,768,1024,768,1024,1024,1024,1024,1024,1024,1024,1024,768,1584,4080,4080,4080,4080,4080,4080,4080,4081,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4080,4080,4064,4080,3520,768,768,1024,768,768,1584,4080,4080,4080,4080,4080,4080,3232,768,768,1024,1024,1024,768,768,1025,1328,3794,4080,4080,4080,4080,4080,4080,4081,1600,768,512,512,512,512,512,512,512,512,256,256,256,256,256,4095),
(0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,513,512,769,512,2688,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4080,4080,4080,4080,2960,768,768,768,1024,1024,768,1856,4080,4080,4080,4080,4080,4080,3793,1040,1025,1025,1024,768,1024,1024,1024,1024,1024,1024,1024,1024,768,2960,4064,4080,4081,4081,4080,4080,2947,1024,768,1024,768,768,4080,4080,4080,4080,4080,4080,768,768,1024,1024,1024,768,768,768,768,768,768,768,768,768,1024,1024,1024,768,768,4080,4080,4080,4080,4080,4080,768,1024,1024,1024,768,768,768,1584,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,3520,768,768,768,1024,1024,1024,1024,1024,1024,1024,1024,768,768,768,768,1024,1024,768,1024,769,768,2976,4080,4081,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,3792,1312,768,768,768,768,1024,768,1024,1024,1024,768,1024,1024,1024,768,768,1584,4080,4080,4080,4080,4080,4081,4080,2976,768,768,768,1024,769,1024,1024,1024,1024,1024,1024,1024,1024,768,1584,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,3521,768,769,1024,768,768,1584,4080,4080,4080,4080,4080,4080,3232,768,768,1024,1024,1024,1024,1024,768,768,2688,4080,4080,4080,4080,4080,4080,4080,3248,512,769,512,512,512,512,512,512,512,256,256,256,256,256,4095),
(0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,514,768,2144,3793,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4080,4080,4065,2416,1040,768,768,1024,768,1024,768,3233,4081,4080,4080,4080,4080,4081,2962,768,768,768,1025,768,1024,1024,1024,1024,1024,1024,1024,1024,768,1856,4082,4080,4080,4080,4080,4080,3808,784,768,1024,769,768,4080,4080,4080,4080,4080,4080,768,1024,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,768,1024,768,768,768,768,4080,4080,4081,4080,4080,4080,768,1024,769,1024,768,768,768,1600,4081,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,3521,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,512,1040,2689,4081,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,3232,1584,768,1025,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,768,1024,768,1024,3778,4080,4080,4080,4080,4080,4082,1584,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,769,768,768,1584,4081,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,3777,768,1025,1024,768,768,1584,4081,4080,4080,4080,4080,4080,3233,768,769,768,768,1024,768,768,769,768,768,3507,4082,4080,4080,4081,4080,4080,4065,2144,512,769,512,512,512,512,512,256,256,256,256,256,256,4095),
(0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,768,768,512,1040,2688,4065,4080,4080,4080,4080,4080,4080,4080,4080,4064,4065,4081,3233,1856,768,768,1024,1024,768,768,768,1312,3794,4080,4064,4080,4080,4080,4065,1856,768,768,768,1024,768,1024,1024,1024,1024,1024,1024,1024,1024,769,1040,3505,4080,4080,4080,4080,4080,4081,2144,768,1024,1024,768,4080,4080,4080,4064,4081,4081,768,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,768,1024,768,768,4065,4080,4081,4080,4080,4081,768,768,1024,1024,1024,768,768,1584,4066,4080,4081,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4080,3777,768,768,1024,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,512,768,2144,3521,4082,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4065,2688,1040,768,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,768,1024,2945,4080,4081,4080,4080,4080,3520,1040,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,768,768,768,1584,4065,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4080,4080,4064,4080,3520,768,768,1024,1024,768,1584,4082,4080,4080,4080,4080,4080,3233,768,768,768,1024,768,768,768,768,768,768,1872,4065,4080,4080,4080,4080,4064,4081,3793,800,256,512,512,512,512,512,256,256,256,256,256,256,4095),
(0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,768,768,512,1056,2416,2960,4064,4064,4080,4081,4081,3792,3248,2960,768,768,768,768,768,768,1024,1025,1024,1024,2144,4066,4080,4080,4080,4064,4066,3779,1040,768,768,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,768,2960,4065,4080,4080,4080,4080,4080,3504,1024,768,1024,768,4080,4080,4080,4080,4081,4048,1040,768,1024,1025,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,768,768,1297,4052,4080,4080,4080,4081,4049,1296,768,768,769,1024,768,1024,1856,4065,4080,4081,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4081,3506,1040,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,769,768,1040,2144,3504,4064,4080,4080,4080,4080,4080,4080,4064,3521,2416,1312,768,768,1024,1024,768,768,768,768,768,768,768,768,768,1024,768,768,1024,768,1024,768,1840,4080,4080,4080,4081,4066,2960,768,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,768,768,1024,1856,4049,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4080,4081,4064,3504,1040,768,1024,1024,1024,1856,4049,4080,4080,4080,4081,4065,3232,1040,768,768,1024,1025,768,768,1024,768,768,768,3235,4082,4064,4080,4080,4080,4080,3808,2432,784,512,512,512,512,512,256,256,256,256,256,256,4095),
(0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,768,512,512,768,512,512,768,768,768,768,768,768,768,768,768,768,770,768,768,768,1024,1025,1024,1024,768,1025,1025,1024,768,768,768,768,1024,1024,768,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1025,768,1024,1024,768,768,768,768,768,768,768,1024,1024,769,1024,768,1024,768,768,1040,769,1024,1024,768,768,768,768,768,768,768,768,768,1024,768,768,1024,768,768,512,1040,768,768,768,1024,1040,513,1024,1024,1024,1024,1024,1025,768,1296,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,512,769,1024,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,769,768,768,768,768,1856,2145,2145,2145,2145,1873,784,768,768,768,1025,1025,768,768,1024,768,768,768,768,768,768,768,768,768,768,768,1024,768,1024,768,1024,768,768,768,768,768,1024,768,1025,768,768,768,768,768,768,768,768,1024,768,1024,1024,768,512,1040,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,768,768,768,1024,1040,768,1024,1024,1024,768,768,1040,768,768,768,768,768,1040,512,1025,1024,1024,768,1024,768,768,768,768,512,768,512,768,768,768,512,512,768,513,513,512,512,512,512,256,256,256,256,256,256,256,4095),
(0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,768,768,512,768,768,512,769,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,768,1024,1024,768,1024,1024,768,1024,768,768,1025,768,768,768,1024,1025,768,768,768,768,768,768,768,768,768,1024,1024,768,768,1024,768,768,768,1024,1024,1024,768,1024,1025,768,768,1025,768,768,1025,768,768,1024,768,768,768,768,768,768,768,768,1024,1024,1024,1024,768,1024,1025,768,768,1024,768,768,1024,1025,1024,768,1024,768,768,1025,768,768,768,1025,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,769,769,768,768,512,768,768,512,768,768,769,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,768,768,768,768,1024,768,768,768,1024,768,768,768,768,768,768,768,768,768,1024,768,768,1024,1024,768,1024,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,1025,768,768,1024,1024,768,1024,1024,1024,768,768,1025,1025,768,768,1024,768,1025,768,768,768,768,768,768,768,512,768,512,769,512,512,768,512,512,512,256,512,512,512,512,512,256,256,256,256,256,256,256,4095),
(0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,768,512,512,512,512,512,768,512,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1025,768,768,768,768,1024,768,768,1024,1024,1024,768,768,1024,1024,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,768,768,1024,768,768,768,768,768,768,1024,768,1024,1024,768,1024,768,1024,768,1024,1024,768,768,768,768,768,768,768,768,768,1024,768,768,1024,1024,768,768,1024,1024,768,1024,768,1024,1024,1024,1024,1024,1024,1024,768,768,768,1025,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,769,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,769,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,768,768,768,1025,1024,768,768,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,1024,768,1024,1024,1024,1024,768,1024,1024,1024,1024,768,768,1024,1024,1024,768,1024,768,768,768,768,768,768,768,768,768,768,768,512,768,512,512,512,512,512,512,512,256,513,256,512,512,512,256,256,256,256,256,256,256,256,4095),
(0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,768,512,512,768,768,512,768,512,512,768,768,768,768,768,768,768,768,768,769,768,768,768,768,768,1024,768,768,1024,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,768,768,768,768,768,1024,768,1024,769,768,1024,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,1024,1024,768,1024,768,768,768,768,768,1024,1024,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,1024,768,768,1024,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,512,512,512,768,512,512,512,512,256,512,512,512,512,256,256,256,256,256,256,256,256,4095),
(0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,768,512,512,512,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,768,768,768,1024,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,768,768,769,768,768,1024,768,768,768,768,768,768,768,768,769,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1025,768,1024,768,768,768,1040,768,768,768,1024,768,768,1024,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,512,512,512,512,768,768,512,768,768,768,768,768,768,768,768,768,768,512,512,768,768,512,769,768,768,768,768,768,768,768,768,768,768,768,768,769,768,768,768,768,768,769,768,768,769,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,769,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,1024,768,768,768,1024,768,1024,768,768,768,768,768,768,769,768,768,768,768,768,768,768,768,768,768,768,768,768,512,512,768,512,512,512,512,512,513,513,512,512,256,512,512,512,256,256,256,256,256,256,256,256,4095),
(0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,4095),
(0,0,0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,4095),
(0,0,0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,256,256,4095),
(0,0,0,0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,768,768,512,512,512,512,512,512,512,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,4095),
(0,0,0,0,0,0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,768,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,0,4095),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,0,0,4095),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,0,0,0,4095),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,0,0,0,4095),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,0,0,0,0,0,4095),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,512,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,256,0,0,0,0,0,0,4095)
);

begin

process(clk)
variable Xoff,Yoff:std_logic_vector(31 downto 0);
begin
if (clk 'event and clk = '1') then
	Xoff := Xpxl - topX;
	Yoff := Ypxl - topY;
	if ( (Xpxl > topX) and (Xpxl < topX + 301) and (Ypxl > topY) and (Ypxl < topY + 71) ) then
		if ( sRGB( conv_integer(Yoff) , conv_integer(Xoff) ) = 0 ) then
			drw <= '0';
		else
			drw <= '1';
			RGB <= conv_std_logic_vector(sRGB(conv_integer(Yoff),conv_integer(Xoff)),12);
		end if;
	else
		drw <= '0';
	end if;
end if;
end process;
end;