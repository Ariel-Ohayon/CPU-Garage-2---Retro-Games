library ieee;
use ieee.std_logic_1164.all;

entity TargetRed is
port(
clk_108:   in  std_logic;
topX,topY: in  std_logic_vector(31 downto 0);
Xpxl,Ypxl: in  std_logic_vector(31 downto 0);
RGB:		  out std_logic_vector(11 downto 0);
drw:		  out std_logic);
end;

architecture one of TargetRed is

component drawTargetRed
port(
clk: in std_logic;
Xpxl,Ypxl: in std_logic_vector(31 downto 0);
topX,topY: in std_logic_vector(31 downto 0);
RGB: out std_logic_vector(11 downto 0);
drw: out std_logic);
end component;

begin
U1: drawTargetRed port map (clk_108,Xpxl,Ypxl,topX,topY,RGB,drw);
end;

-- drawTargetRed
library ieee;
use ieee.std_Logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_Logic_arith.all;

entity drawTargetRed is
port(
clk: in std_logic;
Xpxl,Ypxl: in std_logic_vector(31 downto 0);
topX,topY: in std_logic_vector(31 downto 0);
RGB: out std_logic_vector(11 downto 0);
drw: out std_logic);
end;

architecture one of drawTargetRed is
type mat is array (0 to 164, 0 to 109) of integer range 0 to 4095;
signal sRGB: mat :=
(
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,844,844,844,844,844,844,844,844,844,844,844,844,0,0,0,0,0,0,0,0,844,844,844,844,844,844,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,2577,0,0,0,0,0,0,0,256,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,2577,0,0,0,0,0,0,0,256,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,256,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,256,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,256,0,0,0,0,0,0,0,1280,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,1793,0,0,0,0,1536,1536,1536,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,1793,0,0,0,0,1536,1536,1536,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,1793,0,0,0,0,1536,1536,1536,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,1536,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,1536,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1793,3602,3602,3090,1280,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3602,3602,3602,3602,3602,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0)
);

begin

process(clk)
variable Xoff,Yoff:std_logic_vector(31 downto 0);
begin
if (clk 'event and clk = '1') then
	Xoff := Xpxl - topX;
	Yoff := Ypxl - topY;
	if ( (Xpxl > topX) and (Xpxl < topX + 109) and (Ypxl > topY) and (Ypxl < topY + 164) ) then
		if ( sRGB( conv_integer(Yoff) , conv_integer(Xoff) ) = 0 ) then
			drw <= '0';
		else
			drw <= '1';
			RGB <= conv_std_logic_vector(sRGB(conv_integer(Yoff),conv_integer(Xoff)),12);
		end if;
	else
		drw <= '0';
	end if;
end if;
end process;
end;