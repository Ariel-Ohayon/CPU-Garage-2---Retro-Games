library ieee;
use ieee.std_logic_1164.all;

entity PriorityMux is
port(
P1,P2: 	 in  std_logic_vector(2 downto 0);
in1,in2:  in  std_logic;
l1,l2,l3: out std_logic;
l4,l5,l6: out std_logic);
end;

architecture one of PriorityMux is
signal P: std_logic_vector(5 downto 0);
begin
end;